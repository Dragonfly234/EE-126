library ieee;
use ieee.std_logic_1164.all;


entity MUX64_TB is
end MUX64_TB;

architecture MUX64_TB of MUX64_TB is
 component MUX64
  port(
    in0    : in STD_LOGIC_VECTOR(63 downto 0); 
    in1    : in STD_LOGIC_VECTOR(63 downto 0); 
    sel    : in STD_LOGIC;
    output : out STD_LOGIC_VECTOR(63 downto 0)
);
end component;

signal in0 : STD_LOGIC_VECTOR(63 downto 0):= "0000000000000000000000000000000000000000000000000000000000000000";
signal in1 : STD_LOGIC_VECTOR(63 downto 0):= "0000000000000000000000000000000000000000000000000000000000000000"; 
signal sel:  std_logic:='0';
signal output : STD_LOGIC_VECTOR(63 downto 0);


begin 
   uut: MUX64 port map(
               in0 => in0,
               in1 => in1, 
               output => output,
               sel =>sel
                );


stim_process: process
begin 
  in0 <="0000000000000000000000000000000000000000000000000000000000000000";
  in1 <="1111000000000000000000000000000000000000000000000000000000000000";
  sel<= '1';
  wait for 50 ns;

  in0 <="0000000000000000000000000000000000000000000000000000000000000000";
  in1 <="1010000000000000000000000000000000000000000000000000000000000000";
  sel<= '1';
  wait for 50 ns;

  in0 <="0110000000000000000000000000000000000000000000000000000000000000";
  in1 <="1010000000000000000000000000000000000000000000000000000000000000";
  sel<= '0';
  wait for 50 ns;

  in0 <="1001000000000000000000000000000000000000000000000000000000000000";
  in1 <="0101000000000000000000000000000000000000000000000000000000000000";
  sel<= '0';
  wait ;
end process;
END;
